`timescale 1s/1ms

program test_system_error();

function void main();
    $error;
endfunction : main

initial main();
endprogram : test_system_error
