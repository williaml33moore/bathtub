/*
MIT License

Copyright (c) 2023 Everactive

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in all
copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
SOFTWARE.
*/

`include "bathtub_macros.sv"

// ===================================================================
package bathtub_pkg;
// ===================================================================

	// Main entry point
	`include "bathtub_pkg/bathtub.svh"

	// Resources for step definitions
	`include "bathtub_pkg/step_definition_interface.svh"
	`include "bathtub_pkg/step_static_attributes_interface.svh"
	`include "bathtub_pkg/step_attributes_interface.svh"
	`include "bathtub_pkg/step_nature.svh"
	`include "bathtub_pkg/step_parameters.svh"
	`include "bathtub_pkg/feature_sequence_interface.svh"
	`include "bathtub_pkg/scenario_sequence_interface.svh"

endpackage : bathtub_pkg
