`timescale 1s/1ms

program test_system_fatal();

function void main();
    $fatal;
endfunction : main

initial main();
endprogram : test_system_fatal
